/*************************************************************************************************************
--    Система        : 
--    Разработчик    : 
--    Автор          : Гусев Игорь
--
--    Назначение     : Ram
--------------------------------------------------------------------------------------------------------------
--    Примечание     : 
*************************************************************************************************************/
module ew_ram_r_w_s_dff(
    clk,
    rst_n,
    cs_n,
    wr_n,
    rd_addr,
    wr_addr,
    data_in, 
    data_out
    );

    //----------------------------------------------------------------------//
    // external parameters                                                  //
    //----------------------------------------------------------------------//
    parameter integer DATA_WIDTH    = 32;
    parameter integer RAM_DEPTH     = 8;
    parameter RST_MODE              = 0;
    //----------------------------------------------------------------------//
    // internal parameters                                                  //
    //----------------------------------------------------------------------//
    localparam integer ADDR_WIDTH   = $clog2(RAM_DEPTH);
    //----------------------------------------------------------------------//
    // external signals                                                     //
    //----------------------------------------------------------------------//
    input                           clk;            // входной синхросигнал
    input                           rst_n;          // сигнал сброса
    input                           cs_n;           // подтверждения операции
    input                           wr_n;           // разрешения записи
    input   [ADDR_WIDTH - 1 : 0]    rd_addr;        // шина адреса чтения
    input   [ADDR_WIDTH - 1 : 0]    wr_addr;        // шина адреса записи
    input   [DATA_WIDTH - 1 : 0]    data_in;        // входная шина данных
    output  [DATA_WIDTH - 1 : 0]    data_out;       // выходная шина данных

    //----------------------------------------------------------------------//
    // registers                                                            //
    //----------------------------------------------------------------------//
    reg     [DATA_WIDTH - 1 : 0]    mem [0 : RAM_DEPTH - 1];  // память
    //----------------------------------------------------------------------//
    // assigns                                                              //
    //----------------------------------------------------------------------//
    assign data_out = mem[rd_addr];
    //----------------------------------------------------------------------//
    // logic                                                                //
    //----------------------------------------------------------------------//
    //`ifdef SYNC_MODE_INIT_MEM
    generate 
    if (RST_MODE == 1)
        begin
            always @(posedge clk)
                begin
                    if (~rst_n)  // наивысший приоритет сброс по отрицательному фронту 
                        begin
                            for(int i = 0; i < RAM_DEPTH; i++)
                                mem[i] <= {DATA_WIDTH{1'b0}};
                        end
                    else
                        if (~cs_n &&  ~wr_n)
                            begin
                                mem[wr_addr] <= data_in;
                            end
                end        
        end
    else if (RST_MODE == 0)
        begin
            always @(posedge clk or negedge rst_n)
                begin
                    if (~rst_n)  // наивысший приоритет сброс по отрицательному фронту 
                        begin
                            for(int i = 0; i < RAM_DEPTH; i++)
                                mem[i] <= {DATA_WIDTH{1'b0}};
                        end
                    else
                        if (~cs_n &&  ~wr_n)
                            begin
                                mem[wr_addr] <= data_in;
                            end
                end
        end
    endgenerate

endmodule