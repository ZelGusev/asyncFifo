/*************************************************************************************************************
--    Система        : 
--    Разработчик    : 
--    Автор          : Гусев Игорь
--
--    Назначение     : Управление флагами
--------------------------------------------------------------------------------------------------------------
--    Примечание     : 
*************************************************************************************************************/

module flag(
    clk,
    rst_n,
    data_dm,
    data_dl,
    empty,
    almost_empty,
    half_full,
    almost_full,
    full
    );
    //----------------------------------------------------------------------//
    // external parameters                                                  //
    //----------------------------------------------------------------------//
    parameter integer DATA_WIDTH    = 4;        // ширина шинны данных
    parameter integer RAM_DEPTH     = 8;        // буфер количества слов
    parameter integer AE_LVL        = 2;        // almost empty num word    for write operation
    parameter integer AF_LVL        = 2;        // almost full num word     for write operation
    //----------------------------------------------------------------------//
    // internal parameters                                                  //
    //----------------------------------------------------------------------//
    //----------------------------------------------------------------------//
    // external signals                                                     //
    //----------------------------------------------------------------------//
    input                           clk;
    input                           rst_n;
    input [DATA_WIDTH - 1 : 0]      data_dm;
    input [DATA_WIDTH - 1 : 0]      data_dl;
    output                          empty;
    output                          almost_empty;
    output                          half_full;
    output                          almost_full;
    output                          full;
    //----------------------------------------------------------------------//
    // registers                                                            //
    //----------------------------------------------------------------------//
    //----------------------------------------------------------------------//
    // wire                                                                 //
    //----------------------------------------------------------------------//
    //----------------------------------------------------------------------//
    // assigns                                                              //
    //----------------------------------------------------------------------//
    assign empty        = (data_dm == data_dl);
    assign full         = ((data_dm - data_dl) == RAM_DEPTH);
    assign almost_empty = ((data_dm - data_dl) <= AE_LVL);
    assign half_full    = ((data_dm - data_dl) >= RAM_DEPTH/2);
    assign almost_full  = ((data_dm - data_dl) >= RAM_DEPTH - AF_LVL);
    //----------------------------------------------------------------------//
    // Component instantiations                                             //
    //----------------------------------------------------------------------//
    //----------------------------------------------------------------------//
    // logic                                                                //
    //----------------------------------------------------------------------//
endmodule
