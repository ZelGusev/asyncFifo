/*************************************************************************************************************
--    Система        : 
--    Разработчик    : 
--    Автор          : Гусев Игорь
--
--    Назначение     : Счетчик Грея
--                      С переводом для бинарного счетчика подходит для использования адресации 
--------------------------------------------------------------------------------------------------------------
--    Примечание     : 
*************************************************************************************************************/

module cnt_gray(
    clk,
    rst_n,
    en,
    // msb,
    data_bin,
    data_o
    );
    //----------------------------------------------------------------------//
    // external parameters                                                  //
    //----------------------------------------------------------------------//
    parameter integer DATA_WIDTH    = 4;        // ширина шинны данных
    //----------------------------------------------------------------------//
    // internal parameters                                                  //
    //----------------------------------------------------------------------//
    //----------------------------------------------------------------------//
    // external signals                                                     //
    //----------------------------------------------------------------------//
    input                           clk;
    input                           rst_n;
    input                           en;
    // output reg                      msb;
    output [DATA_WIDTH - 2 : 0]     data_bin;
    output reg [DATA_WIDTH - 1 : 0] data_o;
    //----------------------------------------------------------------------//
    // registers                                                            //
    //----------------------------------------------------------------------//
    //----------------------------------------------------------------------//
    // wire                                                                 //
    //----------------------------------------------------------------------//
    wire [DATA_WIDTH - 1 : 0]  gnext;
    wire [DATA_WIDTH - 1 : 0]  bnext;
    wire [DATA_WIDTH - 1 : 0]  bin;
    //----------------------------------------------------------------------//
    // assigns                                                              //
    //----------------------------------------------------------------------//
    assign bnext    = bin + en;
    assign data_bin = bin;
    //----------------------------------------------------------------------//
    // Component instantiations                                             //
    //----------------------------------------------------------------------//
    grayencode
    #(
        .DATA_WIDTH(DATA_WIDTH)
    )
    grayencode_next
    (
        .data_i     (bnext),
        .data_o     (gnext)
    );
    graydecode
    #(
        .DATA_WIDTH(DATA_WIDTH)
    )
    graydecode_in
    (
        .data_i     (data_o),
        .data_o     (bin)
    );
    //----------------------------------------------------------------------//
    // logic                                                                //
    //----------------------------------------------------------------------//
    `ifdef SYNC_MODE_INIT_MEM
        always @(posedge clk)
            begin
                if (~rst_n)
                    begin
                        data_o  <= {DATA_WIDTH{1'b0}};
                        // msb     <= 1'b0;
                    end
                else
                    begin
                        data_o  <= gnext;
                        // msb     <= gnext[DATA_WIDTH - 2] ^ gnext[DATA_WIDTH - 1];
                    end
            end
    `else
        always @(posedge clk or negedge rst_n)
            begin
                if (~rst_n)
                    begin
                        data_o  <= {DATA_WIDTH{1'b0}};
                        // msb     <= 1'b0;
                    end
                else
                    begin
                        data_o  <= gnext;
                        // msb     <= gnext[DATA_WIDTH - 2] ^ gnext[DATA_WIDTH - 1];
                    end
            end
    `endif
endmodule
