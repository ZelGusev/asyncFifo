/*************************************************************************************************************
--    Система        : 
--    Разработчик    : 
--    Автор          : Гусев Игорь
--
--    Назначение     : encode Grey
--------------------------------------------------------------------------------------------------------------
--    Примечание     : 
*************************************************************************************************************/

module grayencode(
    data_i,
    data_o
    );
    //----------------------------------------------------------------------//
    // external parameters                                                  //
    //----------------------------------------------------------------------//
    parameter integer DATA_WIDTH    = 4;        // ширина шинны данных
    //----------------------------------------------------------------------//
    // internal parameters                                                  //
    //----------------------------------------------------------------------//
    //----------------------------------------------------------------------//
    // external signals                                                     //
    //----------------------------------------------------------------------//
    input  [DATA_WIDTH - 1 : 0]     data_i;
    output  [DATA_WIDTH - 1 : 0]    data_o;
    //----------------------------------------------------------------------//
    // registers                                                            //
    //----------------------------------------------------------------------//
    //----------------------------------------------------------------------//
    // wire                                                                 //
    //----------------------------------------------------------------------//
    //----------------------------------------------------------------------//
    // assigns                                                              //
    //----------------------------------------------------------------------//
    function [DATA_WIDTH - 1 : 0] code;  // соединение информационных данных с проверочными (0)
        input   bit [DATA_WIDTH - 1 : 0]    data;
        begin
            code = data ^ (data >> 1);
        end
    endfunction
    assign data_o = code(data_i);
    //----------------------------------------------------------------------//
    // Component instantiations                                             //
    //----------------------------------------------------------------------//
    //----------------------------------------------------------------------//
    // logic                                                                //
    //----------------------------------------------------------------------//
endmodule
